/***********************************************************************************
 * Copyright (C) 2023 National Research University of Electronic Technology (MIET),
 * Institute of Microdevices and Control Systems.
 * See LICENSE file for licensing details.
 *
 * This file is a part of miriscv core.
 *
 ***********************************************************************************/
import rv_pkg::XLEN;
import rv_gpr_pkg::GPR_ADDR_W;

module rv_control_unit
(
  input  logic                  clk_i,
  input  logic                  arstn_i,

  input  logic [XLEN-1:0]       boot_addr_i,

  input  logic                  f_stall_req_i,
  input  logic                  d_stall_req_i,
  input  logic                  e_stall_req_i,
  input  logic                  m_stall_req_i,

  input  logic [GPR_ADDR_W-1:0] f_cu_rs1_addr_i,
  input  logic                  f_cu_rs1_req_i,
  input  logic [GPR_ADDR_W-1:0] f_cu_rs2_addr_i,
  input  logic                  f_cu_rs2_req_i,

  input  logic [GPR_ADDR_W-1:0] d_cu_rd_addr_i,
  input  logic                  d_cu_rd_we_i,

  input  logic [GPR_ADDR_W-1:0] e_cu_rd_addr_i,
  input  logic                  e_cu_rd_we_i,

  input  logic                  f_valid_i,
  input  logic                  d_valid_i,
  input  logic                  e_valid_i,
  input  logic                  m_valid_i,

  input  logic                  m_branch_i,
  input  logic                  m_jal_i,
  input  logic                  m_jalr_i,
  input  logic [XLEN-1:0]       m_target_pc_i,
  input  logic [XLEN-1:0]       m_next_pc_i,
  input  logic                  m_prediction_i,
  input  logic                  m_br_j_taken_i,

  output logic                  cu_stall_f_o,
  output logic                  cu_stall_d_o,
  output logic                  cu_stall_e_o,
  output logic                  cu_stall_m_o,

  output logic                  cu_kill_f_o,
  output logic                  cu_kill_d_o,
  output logic                  cu_kill_e_o,
  output logic                  cu_kill_m_o,

  output logic [XLEN-1:0]       cu_force_pc_o,
  output logic                  cu_force_f_o
);


  ////////////////////////
  // Local declarations //
  ////////////////////////

  logic [1:0] boot_addr_load_ff;
  logic       cu_boot_addr_load_en;
  logic       cu_mispredict;

  logic       e_raw_hazard_rs1;
  logic       e_raw_hazard_rs2;
  logic       e_raw_hazard;

  logic       m_raw_hazard_rs1;
  logic       m_raw_hazard_rs2;
  logic       m_raw_hazard;


  //////////////////////
  // Pipeline control //
  //////////////////////

  always_ff @(posedge clk_i or negedge arstn_i) begin
    if(~arstn_i) begin
      boot_addr_load_ff <= 2'b00;
    end
    else begin
      boot_addr_load_ff <= {boot_addr_load_ff[0], 1'b1};
    end
  end

  assign cu_boot_addr_load_en = ~boot_addr_load_ff[1];


  assign e_raw_hazard_rs1 = f_cu_rs1_req_i & f_valid_i
                          & d_cu_rd_we_i   & d_valid_i
                          & (f_cu_rs1_addr_i == d_cu_rd_addr_i)
                          & (d_cu_rd_addr_i != '0); // No hazards for x0

  assign e_raw_hazard_rs2 = f_cu_rs2_req_i & f_valid_i
                          & d_cu_rd_we_i   & d_valid_i
                          & (f_cu_rs2_addr_i == d_cu_rd_addr_i)
                          & (d_cu_rd_addr_i != '0); // No hazards for x0


  assign e_raw_hazard = e_raw_hazard_rs1
                      | e_raw_hazard_rs2;

  assign m_raw_hazard_rs1 = f_cu_rs1_req_i & f_valid_i
                          & e_cu_rd_we_i & e_valid_i
                          & (f_cu_rs1_addr_i == e_cu_rd_addr_i)
                          & (e_cu_rd_addr_i != '0); // No hazards for x0

  assign m_raw_hazard_rs2 = f_cu_rs2_req_i & f_valid_i
                          & e_cu_rd_we_i & e_valid_i
                          & (f_cu_rs2_addr_i == e_cu_rd_addr_i)
                          & (e_cu_rd_addr_i != '0); // No hazards for x0

  assign m_raw_hazard = m_raw_hazard_rs1
                      | m_raw_hazard_rs2;


  assign cu_stall_f_o = m_stall_req_i | e_stall_req_i | d_stall_req_i | e_raw_hazard | m_raw_hazard;
  assign cu_stall_d_o = m_stall_req_i | e_stall_req_i | d_stall_req_i;
  assign cu_stall_e_o = m_stall_req_i | e_stall_req_i;
  assign cu_stall_m_o = m_stall_req_i;


  assign cu_mispredict = m_valid_i & (m_prediction_i ^ m_br_j_taken_i) ;

  assign cu_kill_f_o = cu_mispredict;
  assign cu_kill_d_o = cu_mispredict;
  assign cu_kill_e_o = cu_mispredict;
  assign cu_kill_m_o = cu_mispredict;


  assign cu_force_pc_o = cu_boot_addr_load_en ? boot_addr_i
                                              : m_br_j_taken_i ? m_target_pc_i
                                                               : m_next_pc_i;

  assign cu_force_f_o = cu_boot_addr_load_en | cu_mispredict;

endmodule