/***********************************************************************************
 * Copyright (C) 2023 National Research University of Electronic Technology (MIET),
 * Institute of Microdevices and Control Systems.
 * See LICENSE file for licensing details.
 *
 * This file is a part of miriscv core.
 *
 ***********************************************************************************/

package  rv_gpr_pkg;

  parameter     GPR_ADDR_W  = 5;    // GPR address width

endpackage :  rv_gpr_pkg